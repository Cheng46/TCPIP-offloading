
module igmp_client(
    input wire      i_sys_clk,
    input wire      i_rstn,

    
);

endmodule